



`timescale 1ns/1ps

module tb_udp_parser;

    localparam DEPTH = 31;

    // Input signals
    logic clock;
    logic reset;
    logic [255:0] a_data_i;
    logic a_valid_i;
    logic out_ready;
    // Output signals
    logic a_ready_o;
    logic b_ready_i;
    logic [31:0] b_data_o;
    logic b_valid_o;
    
    udp_parser dut
    (
        .clock          (clock),
        .reset          (reset),
        .a_data_i       (a_data_i),
        .a_valid_i      (a_valid_i),
        .b_ready_i      (b_ready_i),
        .b_data_o       (b_data_o),
        .b_valid_o      (b_valid_o)
    );
        
    task generate_sequence;
    begin
        $display("Starting simple input sequence");
        @(posedge clock) a_valid_i<= 1'b1;
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{32'b10},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        @(posedge clock) a_data_i <= {{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1},{{DEPTH{1'b0}},1'b1}};
        $display("Simple input sequence done");
    end
    endtask

    // Clock generation
    always begin
        #5 clock = ~clock;
    end

    // Test stimulus generation
    initial begin
        // Initialize inputs
        clock = 0;
        reset = 1'b1;
        a_valid_i = 1'b0;
        b_ready_i = 1'b1;
        a_data_i = 0;

        // Apply reset
        #10 reset = 0;
        generate_sequence();
        repeat(10) @(posedge clock);
        $finish;
    end
endmodule


       